/*
*Author : Revanth Sai Nandamuri
*Portfolio : https://revanthnandamuri1341b0.github.io/
*Date of update : 24 January 2022
*Project name : 
*Domain : 
*Description : Pre-Defined Sequencer
*File Name : sequencer.sv
*File ID : 644159
*Modified by : #your name#
*/
typedef uvm_sequencer #(packet) sequencer;